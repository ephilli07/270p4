`timescale 1ns/1ns

module TestBenchFullAdder( 

);


FullAdder testFullAdder(); 

initial begin 
    
end

endmodule