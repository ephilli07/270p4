// File Name: CombCalc.v
module  CombCalc(
	input [2:0] OP,
	input signed [3:0] A, B,
	output signed [3:0] R,
	output ovf
);

	wire signed [3:0] X, Y;
	wire c0;

// Prefix Circuit


// Instantiate a 4-bit Adder/Subtractor

endmodule //  CombCalc